----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:05:46 09/30/2016 
-- Design Name: 
-- Module Name:    count1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity count1 is
    Port ( sw : in  STD_LOGIC_VECTOR (7 downto 0);
           res : out  STD_LOGIC_VECTOR (3 downto 0));
end count1;

architecture Behavioral of count1 is

begin

	PROCESS(sw)
	VARIABLE count1_res : INTEGER;
	BEGIN
			count1_res := 0;
			loop_count1: FOR cpt IN 0 TO 7 LOOP
				if sw(cpt) = '1' then count1_res := count1_res + 1; end if;
			END LOOP loop_count1;
			res <= conv_std_logic_vector(count1_res, 4);
	END PROCESS; 


end Behavioral;

